

module ether_tx(
	clk_50M,
	tx_en,
	tx_d
);

	input clk_50M;
	output tx_en;
	output [1:0] tx_d;

endmodule
