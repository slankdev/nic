

module ether_rx(
	clk_50M,
	rx_dv,
	rx_d
);

	input clk_50M;
	input rx_dv;
	input [1:0] rx_d;

endmodule
